magic
tech sky130B
magscale 1 2
timestamp 1686891616
<< nwell >>
rect 7000 6462 8090 10722
rect 7000 6438 8124 6462
rect 7000 4058 7056 6438
rect 7144 4126 7202 4184
rect 8024 4178 8124 6438
rect 7996 4100 8454 4178
rect 8466 4122 8540 4200
rect 8024 4060 8124 4100
<< pwell >>
rect 6330 9196 6800 9986
rect 8940 7000 10120 9586
rect 6980 3360 7070 3400
rect 6980 3238 7022 3360
rect 6980 3218 7070 3238
rect 6980 2640 7022 3218
rect 7460 2810 7622 3168
rect 7036 2664 7116 2730
rect 9100 2440 9160 6704
rect 9920 4000 10120 6704
rect 6400 2422 7000 2440
rect 8042 2422 8070 2440
rect 6400 2420 7036 2422
rect 6992 2400 7036 2420
rect 8042 2400 8078 2422
rect 6992 2388 7106 2400
rect 8024 2388 8078 2400
rect 6992 2384 7126 2388
rect 6450 2070 6504 2210
rect 6450 2066 6500 2070
rect 6450 70 6544 2066
rect 6500 66 6544 70
rect 6956 36 7166 2384
rect 7866 210 7886 2210
rect 7948 2198 8078 2388
rect 7900 1864 7946 1898
rect 7514 122 7576 190
rect 7954 96 8078 2198
rect 9536 122 9594 186
rect 7900 48 8078 96
rect 6992 0 7118 36
rect 7954 0 8078 48
rect 9930 46 9990 4000
rect 9140 0 9990 46
<< psubdiff >>
rect 6956 36 7166 2384
<< poly >>
rect 8466 4122 8540 4200
rect 7514 122 7576 190
rect 9536 122 9594 186
<< locali >>
rect 5000 10912 10120 10972
rect 5000 10712 5300 10912
rect 9954 10712 10120 10912
rect 5000 10652 10120 10712
rect 5000 10200 8148 10652
rect 5000 9950 6800 10000
rect 5000 9800 5540 9950
rect 5000 1000 5064 9800
rect 5264 4826 5540 9800
rect 6278 9160 6800 9950
rect 6260 9150 6800 9160
rect 5264 1000 5566 4826
rect 5000 848 5566 1000
rect 6260 4070 6400 9150
rect 6758 4070 6800 9150
rect 6260 4000 6800 4070
rect 7000 6368 8148 10200
rect 8858 7000 10120 10652
rect 7000 4070 7056 6368
rect 8024 4070 8124 6368
rect 8858 4070 8940 7000
rect 7000 4000 8940 4070
rect 9100 6644 10120 6704
rect 6260 848 6330 4000
rect 6980 3390 8100 3400
rect 6980 3350 7200 3390
rect 7878 3350 8100 3390
rect 6980 3332 8100 3350
rect 6980 2640 7070 3332
rect 8026 2640 8100 3332
rect 6980 2636 7460 2640
rect 7620 2636 8100 2640
rect 6980 2630 8100 2636
rect 6980 2590 7036 2630
rect 8042 2590 8100 2630
rect 6980 2580 8100 2590
rect 9100 3200 9210 6644
rect 9100 3164 9180 3200
rect 9100 2440 9186 3164
rect 5000 790 6330 848
rect 6390 2436 9186 2440
rect 6390 2374 9176 2436
rect 6390 400 6490 2374
rect 5000 70 6490 400
rect 6956 70 7166 2374
rect 7866 2370 9176 2374
rect 7932 1898 9176 2370
rect 7900 1864 9176 1898
rect 7932 96 9176 1864
rect 7900 70 9176 96
rect 9920 70 10120 6644
rect 5000 0 10120 70
rect 5000 -200 5300 0
rect 9954 -200 10120 0
rect 5000 -250 10120 -200
<< viali >>
rect 5300 10712 9954 10912
rect 5064 1000 5264 9800
rect 7200 3350 7878 3390
rect 7036 2590 8042 2630
rect 5300 -200 9954 0
<< metal1 >>
rect 9384 11200 9394 11400
rect 9594 11200 9604 11400
rect 5000 10912 10120 10972
rect 5000 10712 5300 10912
rect 9954 10712 10120 10912
rect 5000 10652 10120 10712
rect 5000 9800 5320 10000
rect 5000 1000 5064 9800
rect 5264 1000 5320 9800
rect 5628 9388 5834 10652
rect 6026 9388 6634 9820
rect 6496 8598 6634 9388
rect 7460 6220 7620 10652
rect 8166 10504 8216 10652
rect 6496 2800 6634 4598
rect 7080 4218 7190 6220
rect 7402 4218 7676 6220
rect 7888 4218 7998 6220
rect 8166 4218 8268 10504
rect 7080 4184 7144 4218
rect 7080 4126 7878 4184
rect 7934 4178 7998 4218
rect 8350 4178 8400 10544
rect 8464 4218 8474 10504
rect 8532 4218 8542 10504
rect 8606 4178 8656 10544
rect 8790 10504 8840 10652
rect 8738 4218 8840 10504
rect 9412 6532 9462 6544
rect 9670 6532 9720 6544
rect 9370 6526 9500 6532
rect 9630 6526 9760 6532
rect 7080 2990 7144 4126
rect 7934 4100 8732 4178
rect 7188 3390 7890 3396
rect 7188 3350 7200 3390
rect 7878 3350 7890 3390
rect 7188 3344 7890 3350
rect 7460 3308 7620 3344
rect 7080 2810 7190 2990
rect 7230 2814 7360 3200
rect 6496 2600 6948 2800
rect 7230 2732 7260 2814
rect 7340 2732 7360 2814
rect 7402 2810 7500 3168
rect 7590 2810 7676 3168
rect 7718 2820 7848 3200
rect 7934 2990 7998 4100
rect 7718 2772 7740 2820
rect 7730 2738 7740 2772
rect 7820 2772 7848 2820
rect 7888 2810 7998 2990
rect 7820 2738 7830 2772
rect 5000 790 5320 1000
rect 5662 956 6164 1388
rect 6450 70 6544 2210
rect 6630 178 6760 2242
rect 6854 2210 6948 2600
rect 7024 2630 8054 2636
rect 7024 2590 7036 2630
rect 8042 2590 8054 2630
rect 7024 2584 8054 2590
rect 7350 2244 7480 2248
rect 7350 2242 7440 2244
rect 7608 2242 7738 2248
rect 6848 210 6948 2210
rect 7200 290 7262 2210
rect 7200 230 7220 290
rect 7280 230 7290 290
rect 7200 210 7262 230
rect 6854 178 6948 210
rect 7390 178 7440 2242
rect 7490 222 7500 2210
rect 7590 222 7600 2210
rect 7648 178 7698 2242
rect 7824 290 7886 2210
rect 7796 230 7806 290
rect 7866 230 7886 290
rect 7824 210 7886 230
rect 9240 280 9330 6494
rect 9240 220 9260 280
rect 9320 220 9330 280
rect 9240 210 9330 220
rect 9412 178 9462 6526
rect 9526 210 9536 6496
rect 9594 210 9604 6496
rect 9670 178 9720 6526
rect 9800 210 9890 6494
rect 6596 110 9794 178
rect 9852 70 9890 210
rect 5000 40 10120 70
rect 5000 0 7220 40
rect 7280 0 7806 40
rect 7866 0 9260 40
rect 9320 0 10120 40
rect 5000 -200 5300 0
rect 9954 -200 10120 0
rect 5000 -250 10120 -200
rect 6906 -600 6916 -400
rect 7116 -600 7126 -400
rect 7954 -600 7964 -400
rect 8164 -600 8174 -400
<< via1 >>
rect 9394 11200 9594 11400
rect 8474 4218 8532 10504
rect 7260 2732 7340 2814
rect 7500 2810 7590 3168
rect 7740 2738 7820 2820
rect 7220 230 7280 290
rect 7500 222 7590 2210
rect 7806 230 7866 290
rect 9260 220 9320 280
rect 9536 210 9594 6496
rect 7220 0 7280 40
rect 7806 0 7866 40
rect 9260 0 9320 40
rect 7220 -20 7280 0
rect 7806 -20 7866 0
rect 9260 -20 9320 0
rect 6916 -600 7116 -400
rect 7964 -600 8164 -400
<< metal2 >>
rect 9394 11400 9594 11410
rect 9394 10514 9594 11200
rect 8474 10504 9594 10514
rect 8532 6496 9594 10504
rect 8532 4218 9536 6496
rect 8474 4208 9536 4218
rect 7500 3168 7590 3178
rect 6916 2814 7340 2824
rect 6916 2732 7260 2814
rect 6916 2722 7340 2732
rect 6916 -400 7116 2722
rect 7500 2210 7590 2810
rect 7740 2820 8164 2830
rect 7820 2738 8164 2820
rect 7740 2728 8164 2738
rect 7220 290 7280 300
rect 7220 40 7280 230
rect 7500 212 7590 222
rect 7806 290 7866 300
rect 7220 -30 7280 -20
rect 7806 40 7866 230
rect 7806 -30 7866 -20
rect 6916 -610 7116 -600
rect 7964 -400 8164 2728
rect 9260 280 9320 290
rect 9260 40 9320 220
rect 9536 200 9594 210
rect 9260 -30 9320 -20
rect 7964 -610 8164 -600
use sky130_fd_pr__nfet_01v8_34YWRA  xm1
timestamp 1685705005
transform 1 0 7296 0 1 2989
box -296 -389 296 389
use sky130_fd_pr__nfet_01v8_34YWRA  xm2
timestamp 1685705005
transform 1 0 7782 0 1 2989
box -296 -389 296 389
use sky130_fd_pr__pfet_01v8_GGAEPD  xm3
timestamp 1685705005
transform 1 0 7296 0 1 5219
box -296 -1219 296 1219
use sky130_fd_pr__pfet_01v8_GGAEPD  xm4
timestamp 1685705005
transform 1 0 7782 0 1 5219
box -296 -1219 296 1219
use sky130_fd_pr__nfet_01v8_EF4BLE  xm5
timestamp 1685705005
transform 1 0 7543 0 1 1210
box -425 -1210 425 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  xm6
timestamp 1685705005
transform 1 0 6696 0 1 1210
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_RLGYC7  xm7
timestamp 1685705005
transform 1 0 8503 0 1 7361
box -425 -3361 425 3361
use sky130_fd_pr__nfet_01v8_6WGMFU  xm8
timestamp 1685705005
transform 1 0 9565 0 1 3352
box -425 -3352 425 3352
use sky130_fd_pr__res_high_po_0p69_NKSDAM  xR1
timestamp 1685705005
transform 1 0 5731 0 1 5388
box -235 -4598 235 4598
use sky130_fd_pr__res_high_po_0p69_NKSDAM  xR2
timestamp 1685705005
transform 1 0 6095 0 1 5388
box -235 -4598 235 4598
use sky130_fd_pr__res_high_po_0p69_YVB7ZU  xR3
timestamp 1685705005
transform 1 0 6565 0 1 6598
box -235 -2598 235 2598
<< labels >>
flabel metal1 5000 -200 5200 0 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 5000 10712 5200 10912 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel via1 9394 11200 9594 11400 0 FreeSans 256 0 0 0 out2
port 5 nsew
flabel via1 6916 -600 7116 -400 0 FreeSans 256 0 0 0 in1
port 3 nsew
flabel via1 7964 -600 8164 -400 0 FreeSans 256 0 0 0 in2
port 4 nsew
flabel metal1 5064 5202 5264 5402 0 FreeSans 256 0 0 0 vss
<< end >>
