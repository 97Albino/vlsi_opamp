magic
tech sky130B
magscale 1 2
timestamp 1685705005
<< nwell >>
rect -296 -1219 296 1219
<< pmos >>
rect -100 -1000 100 1000
<< pdiff >>
rect -158 988 -100 1000
rect -158 -988 -146 988
rect -112 -988 -100 988
rect -158 -1000 -100 -988
rect 100 988 158 1000
rect 100 -988 112 988
rect 146 -988 158 988
rect 100 -1000 158 -988
<< pdiffc >>
rect -146 -988 -112 988
rect 112 -988 146 988
<< nsubdiff >>
rect -260 1149 -164 1183
rect 164 1149 260 1183
rect -260 1087 -226 1149
rect 226 1087 260 1149
rect -260 -1149 -226 -1087
rect 226 -1149 260 -1087
rect -260 -1183 -164 -1149
rect 164 -1183 260 -1149
<< nsubdiffcont >>
rect -164 1149 164 1183
rect -260 -1087 -226 1087
rect 226 -1087 260 1087
rect -164 -1183 164 -1149
<< poly >>
rect -100 1081 100 1097
rect -100 1047 -84 1081
rect 84 1047 100 1081
rect -100 1000 100 1047
rect -100 -1047 100 -1000
rect -100 -1081 -84 -1047
rect 84 -1081 100 -1047
rect -100 -1097 100 -1081
<< polycont >>
rect -84 1047 84 1081
rect -84 -1081 84 -1047
<< locali >>
rect -260 1149 -164 1183
rect 164 1149 260 1183
rect -260 1087 -226 1149
rect 226 1087 260 1149
rect -100 1047 -84 1081
rect 84 1047 100 1081
rect -146 988 -112 1004
rect -146 -1004 -112 -988
rect 112 988 146 1004
rect 112 -1004 146 -988
rect -100 -1081 -84 -1047
rect 84 -1081 100 -1047
rect -260 -1149 -226 -1087
rect 226 -1149 260 -1087
rect -260 -1183 -164 -1149
rect 164 -1183 260 -1149
<< viali >>
rect -84 1047 84 1081
rect -146 -988 -112 988
rect 112 -988 146 988
rect -84 -1081 84 -1047
<< metal1 >>
rect -96 1081 96 1087
rect -96 1047 -84 1081
rect 84 1047 96 1081
rect -96 1041 96 1047
rect -152 988 -106 1000
rect -152 -988 -146 988
rect -112 -988 -106 988
rect -152 -1000 -106 -988
rect 106 988 152 1000
rect 106 -988 112 988
rect 146 -988 152 988
rect 106 -1000 152 -988
rect -96 -1047 96 -1041
rect -96 -1081 -84 -1047
rect 84 -1081 96 -1047
rect -96 -1087 96 -1081
<< properties >>
string FIXED_BBOX -243 -1166 243 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
