magic
tech sky130B
magscale 1 2
timestamp 1685705005
<< pwell >>
rect -425 -3352 425 3352
<< nmos >>
rect -229 -3142 -29 3142
rect 29 -3142 229 3142
<< ndiff >>
rect -287 3130 -229 3142
rect -287 -3130 -275 3130
rect -241 -3130 -229 3130
rect -287 -3142 -229 -3130
rect -29 3130 29 3142
rect -29 -3130 -17 3130
rect 17 -3130 29 3130
rect -29 -3142 29 -3130
rect 229 3130 287 3142
rect 229 -3130 241 3130
rect 275 -3130 287 3130
rect 229 -3142 287 -3130
<< ndiffc >>
rect -275 -3130 -241 3130
rect -17 -3130 17 3130
rect 241 -3130 275 3130
<< psubdiff >>
rect -389 3282 -293 3316
rect 293 3282 389 3316
rect -389 3220 -355 3282
rect 355 3220 389 3282
rect -389 -3282 -355 -3220
rect 355 -3282 389 -3220
rect -389 -3316 -293 -3282
rect 293 -3316 389 -3282
<< psubdiffcont >>
rect -293 3282 293 3316
rect -389 -3220 -355 3220
rect 355 -3220 389 3220
rect -293 -3316 293 -3282
<< poly >>
rect -229 3214 -29 3230
rect -229 3180 -213 3214
rect -45 3180 -29 3214
rect -229 3142 -29 3180
rect 29 3214 229 3230
rect 29 3180 45 3214
rect 213 3180 229 3214
rect 29 3142 229 3180
rect -229 -3180 -29 -3142
rect -229 -3214 -213 -3180
rect -45 -3214 -29 -3180
rect -229 -3230 -29 -3214
rect 29 -3180 229 -3142
rect 29 -3214 45 -3180
rect 213 -3214 229 -3180
rect 29 -3230 229 -3214
<< polycont >>
rect -213 3180 -45 3214
rect 45 3180 213 3214
rect -213 -3214 -45 -3180
rect 45 -3214 213 -3180
<< locali >>
rect -389 3282 -293 3316
rect 293 3282 389 3316
rect -389 3220 -355 3282
rect 355 3220 389 3282
rect -229 3180 -213 3214
rect -45 3180 -29 3214
rect 29 3180 45 3214
rect 213 3180 229 3214
rect -275 3130 -241 3146
rect -275 -3146 -241 -3130
rect -17 3130 17 3146
rect -17 -3146 17 -3130
rect 241 3130 275 3146
rect 241 -3146 275 -3130
rect -229 -3214 -213 -3180
rect -45 -3214 -29 -3180
rect 29 -3214 45 -3180
rect 213 -3214 229 -3180
rect -389 -3282 -355 -3220
rect 355 -3282 389 -3220
rect -389 -3316 -293 -3282
rect 293 -3316 389 -3282
<< viali >>
rect -213 3180 -45 3214
rect 45 3180 213 3214
rect -275 -3130 -241 3130
rect -17 -3130 17 3130
rect 241 -3130 275 3130
rect -213 -3214 -45 -3180
rect 45 -3214 213 -3180
<< metal1 >>
rect -225 3214 -33 3220
rect -225 3180 -213 3214
rect -45 3180 -33 3214
rect -225 3174 -33 3180
rect 33 3214 225 3220
rect 33 3180 45 3214
rect 213 3180 225 3214
rect 33 3174 225 3180
rect -281 3130 -235 3142
rect -281 -3130 -275 3130
rect -241 -3130 -235 3130
rect -281 -3142 -235 -3130
rect -23 3130 23 3142
rect -23 -3130 -17 3130
rect 17 -3130 23 3130
rect -23 -3142 23 -3130
rect 235 3130 281 3142
rect 235 -3130 241 3130
rect 275 -3130 281 3130
rect 235 -3142 281 -3130
rect -225 -3180 -33 -3174
rect -225 -3214 -213 -3180
rect -45 -3214 -33 -3180
rect -225 -3220 -33 -3214
rect 33 -3180 225 -3174
rect 33 -3214 45 -3180
rect 213 -3214 225 -3180
rect 33 -3220 225 -3214
<< properties >>
string FIXED_BBOX -372 -3299 372 3299
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 31.415 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
