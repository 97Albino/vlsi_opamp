magic
tech sky130B
magscale 1 2
timestamp 1686918407
<< nwell >>
rect -425 -3361 425 3361
<< pmos >>
rect -229 -3142 -29 3142
rect 29 -3142 229 3142
<< pdiff >>
rect -287 3130 -229 3142
rect -287 -3130 -275 3130
rect -241 -3130 -229 3130
rect -287 -3142 -229 -3130
rect -29 3130 29 3142
rect -29 -3130 -17 3130
rect 17 -3130 29 3130
rect -29 -3142 29 -3130
rect 229 3130 287 3142
rect 229 -3130 241 3130
rect 275 -3130 287 3130
rect 229 -3142 287 -3130
<< pdiffc >>
rect -275 -3130 -241 3130
rect -17 -3130 17 3130
rect 241 -3130 275 3130
<< nsubdiff >>
rect -389 3291 -293 3325
rect 293 3291 389 3325
rect -389 3229 -355 3291
rect 355 3229 389 3291
rect -389 -3291 -355 -3229
rect 355 -3291 389 -3229
rect -389 -3325 -293 -3291
rect 293 -3325 389 -3291
<< nsubdiffcont >>
rect -293 3291 293 3325
rect -389 -3229 -355 3229
rect 355 -3229 389 3229
rect -293 -3325 293 -3291
<< poly >>
rect -229 3223 -29 3239
rect -229 3189 -213 3223
rect -45 3189 -29 3223
rect -229 3142 -29 3189
rect 29 3223 229 3239
rect 29 3189 45 3223
rect 213 3189 229 3223
rect 29 3142 229 3189
rect -229 -3189 -29 -3142
rect -229 -3223 -213 -3189
rect -45 -3223 -29 -3189
rect -229 -3239 -29 -3223
rect 29 -3189 229 -3142
rect 29 -3223 45 -3189
rect 213 -3223 229 -3189
rect 29 -3239 229 -3223
<< polycont >>
rect -213 3189 -45 3223
rect 45 3189 213 3223
rect -213 -3223 -45 -3189
rect 45 -3223 213 -3189
<< locali >>
rect -389 3291 -293 3325
rect 293 3291 389 3325
rect -389 3229 -355 3291
rect 355 3229 389 3291
rect -229 3189 -213 3223
rect -45 3189 -29 3223
rect 29 3189 45 3223
rect 213 3189 229 3223
rect -275 3130 -241 3146
rect -275 -3146 -241 -3130
rect -17 3130 17 3146
rect -17 -3146 17 -3130
rect 241 3130 275 3146
rect 241 -3146 275 -3130
rect -229 -3223 -213 -3189
rect -45 -3223 -29 -3189
rect 29 -3223 45 -3189
rect 213 -3223 229 -3189
rect -389 -3291 -355 -3229
rect 355 -3291 389 -3229
rect -389 -3325 -293 -3291
rect 293 -3325 389 -3291
<< viali >>
rect -213 3189 -45 3223
rect 45 3189 213 3223
rect -275 -3130 -241 3130
rect -17 -3130 17 3130
rect 241 -3130 275 3130
rect -213 -3223 -45 -3189
rect 45 -3223 213 -3189
<< metal1 >>
rect -225 3223 -33 3229
rect -225 3189 -213 3223
rect -45 3189 -33 3223
rect -225 3183 -33 3189
rect 33 3223 225 3229
rect 33 3189 45 3223
rect 213 3189 225 3223
rect 33 3183 225 3189
rect -281 3130 -235 3142
rect -281 -3130 -275 3130
rect -241 -3130 -235 3130
rect -281 -3142 -235 -3130
rect -23 3130 23 3142
rect -23 -3130 -17 3130
rect 17 -3130 23 3130
rect -23 -3142 23 -3130
rect 235 3130 281 3142
rect 235 -3130 241 3130
rect 275 -3130 281 3130
rect 235 -3142 281 -3130
rect -225 -3189 -33 -3183
rect -225 -3223 -213 -3189
rect -45 -3223 -33 -3189
rect -225 -3229 -33 -3223
rect 33 -3189 225 -3183
rect 33 -3223 45 -3189
rect 213 -3223 225 -3189
rect 33 -3229 225 -3223
<< properties >>
string FIXED_BBOX -372 -3308 372 3308
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 31.415 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
