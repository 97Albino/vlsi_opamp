.subckt res r0 r1 gnd
r0 r1 gnd sky130_fd_pr__res_high_po_0p69 l=5
.ends
