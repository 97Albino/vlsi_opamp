magic
tech sky130B
magscale 1 2
timestamp 1686928317
<< nwell >>
rect 7300 9446 8288 9922
rect 7300 5592 8324 9446
rect 7300 3256 7368 5592
rect 8668 3322 8726 3400
<< pwell >>
rect 6000 9126 7198 9196
rect 6000 36 6042 9126
rect 6808 7494 7198 9126
rect 7148 3092 7198 7458
rect 7128 3044 9268 3092
rect 6894 2480 7070 2912
rect 7128 2352 7336 3044
rect 8262 2384 9268 3044
rect 7128 2350 7484 2352
rect 7250 36 7484 2350
rect 8194 70 9270 2384
rect 9942 70 9980 214
rect 7292 0 7432 36
rect 8194 0 10080 70
<< psubdiff >>
rect 6000 9126 7198 9196
rect 6000 36 6042 9126
rect 7128 3044 9268 3092
rect 7128 2352 7336 3044
rect 8308 2384 9268 3044
rect 7128 2350 7484 2352
rect 7250 36 7484 2350
rect 8194 70 9270 2384
rect 8194 0 10080 70
<< poly >>
rect 8668 3322 8726 3400
<< locali >>
rect 6000 10120 10080 10182
rect 6000 9920 6260 10120
rect 9880 9920 10080 10120
rect 6000 9852 10080 9920
rect 6000 9300 8324 9852
rect 6000 9126 7198 9196
rect 6000 70 6042 9126
rect 6786 7446 7198 9126
rect 7148 3092 7198 7446
rect 7300 5592 8324 9300
rect 9064 6800 10080 9852
rect 7300 3270 7368 5592
rect 9072 3270 9122 6800
rect 7300 3200 9122 3270
rect 9230 6636 10080 6704
rect 9230 3092 9284 6636
rect 7128 3044 9268 3092
rect 7128 2352 7336 3044
rect 8308 2384 9268 3044
rect 7128 2350 7484 2352
rect 7250 70 7484 2350
rect 8194 70 9270 2384
rect 10026 70 10080 6636
rect 6000 0 10080 70
rect 6000 -200 6260 0
rect 9880 -200 10080 0
rect 6000 -260 10080 -200
<< viali >>
rect 6260 9920 9880 10120
rect 6260 -200 9880 0
<< metal1 >>
rect 9490 10300 9500 10500
rect 9700 10300 9710 10500
rect 6000 10120 10080 10182
rect 6000 9920 6260 10120
rect 9880 9920 10080 10120
rect 6000 9852 10080 9920
rect 6166 8598 6304 9852
rect 6530 8598 7032 9030
rect 6894 6912 7032 8598
rect 7400 3418 7490 5420
rect 7400 3378 7444 3418
rect 7540 3378 7650 5490
rect 7760 5420 7920 9852
rect 8360 9704 8410 9852
rect 8520 9744 8620 9778
rect 8780 9744 8880 9778
rect 7702 3418 7976 5420
rect 7400 3332 7992 3378
rect 8030 3374 8140 5490
rect 8234 3378 8278 5420
rect 8360 3418 8462 9704
rect 8520 3380 8600 9744
rect 8650 3418 8660 9704
rect 8734 3418 8744 9704
rect 8234 3332 8484 3378
rect 8520 3332 8620 3380
rect 8800 3378 8880 9744
rect 8984 9704 9040 9852
rect 8932 3418 9040 9704
rect 8780 3332 8880 3378
rect 6894 2242 7180 2912
rect 7400 2524 7444 3332
rect 7560 2492 7640 2916
rect 7702 2860 7976 2882
rect 7702 2540 7800 2860
rect 7880 2540 7976 2860
rect 7702 2524 7976 2540
rect 8044 2492 8124 2926
rect 8234 2524 8278 3332
rect 7490 2432 7500 2492
rect 7692 2432 7702 2492
rect 7976 2432 7986 2492
rect 8178 2432 8188 2492
rect 6166 166 6668 598
rect 6780 70 6878 2210
rect 6960 178 7180 2242
rect 7518 280 7604 2210
rect 7518 220 7528 280
rect 7588 220 7604 280
rect 7518 210 7604 220
rect 7680 178 7740 2246
rect 7790 210 7800 2210
rect 7880 210 7890 2210
rect 7940 178 8000 2246
rect 8074 280 8160 2210
rect 8074 220 8090 280
rect 8150 220 8160 280
rect 8074 210 8160 220
rect 9328 282 9374 6494
rect 9328 222 9342 282
rect 9402 222 9412 282
rect 9328 210 9374 222
rect 9616 210 9626 6494
rect 9684 210 9694 6494
rect 9890 210 10000 6494
rect 6928 132 9752 178
rect 9942 70 10000 210
rect 6000 60 10080 70
rect 6000 0 7528 60
rect 7588 0 8090 60
rect 8150 0 9342 60
rect 9402 0 10080 60
rect 6000 -200 6260 0
rect 9880 -200 10080 0
rect 6000 -260 10080 -200
rect 7210 -546 7220 -346
rect 7420 -546 7430 -346
rect 8258 -546 8268 -346
rect 8468 -546 8478 -346
<< via1 >>
rect 9500 10300 9700 10500
rect 8660 3418 8734 9704
rect 7800 2540 7880 2860
rect 7500 2432 7692 2492
rect 7986 2432 8178 2492
rect 7528 220 7588 280
rect 7800 210 7880 2210
rect 8090 220 8150 280
rect 9342 222 9402 282
rect 9626 210 9684 6494
rect 7528 0 7588 60
rect 8090 0 8150 60
rect 9342 0 9402 60
rect 7220 -546 7420 -346
rect 8268 -546 8468 -346
<< metal2 >>
rect 9500 10500 9700 10510
rect 9500 9714 9700 10300
rect 8660 9704 9700 9714
rect 8734 6494 9700 9704
rect 8734 3418 9626 6494
rect 7800 2860 7880 2870
rect 7220 2492 7692 2502
rect 7220 2432 7500 2492
rect 7220 2422 7692 2432
rect 7220 -346 7420 2422
rect 7800 2210 7880 2540
rect 7986 2492 8468 2502
rect 8178 2432 8468 2492
rect 7986 2422 8468 2432
rect 7528 280 7588 290
rect 7528 60 7588 220
rect 7800 200 7880 210
rect 8090 280 8150 290
rect 7528 -10 7588 0
rect 8090 60 8150 220
rect 8090 -10 8150 0
rect 7220 -556 7420 -546
rect 8268 -346 8468 2422
rect 8660 520 9626 3418
rect 9342 282 9402 292
rect 9342 60 9402 222
rect 9520 210 9626 520
rect 9684 210 9700 6494
rect 9520 200 9700 210
rect 9342 -10 9402 0
rect 8268 -556 8468 -546
use sky130_fd_pr__nfet_01v8_RXBUCF  sky130_fd_pr__nfet_01v8_RXBUCF_0
timestamp 1686927284
transform 1 0 7596 0 1 2703
box -296 -389 296 389
use sky130_fd_pr__nfet_01v8_RXBUCF  xm2
timestamp 1686927284
transform 1 0 8082 0 1 2703
box -296 -389 296 389
use sky130_fd_pr__pfet_01v8_GGAEPD  xm3
timestamp 1686918407
transform 1 0 7596 0 1 4419
box -296 -1219 296 1219
use sky130_fd_pr__pfet_01v8_GABEPD  xm4
timestamp 1686927284
transform 1 0 8082 0 1 4419
box -296 -1219 296 1219
use sky130_fd_pr__nfet_01v8_EF4BLE  xm5
timestamp 1686918407
transform 1 0 7839 0 1 1210
box -425 -1210 425 1210
use sky130_fd_pr__nfet_01v8_9FXQ3X  xm6
timestamp 1686918407
transform 1 0 7024 0 1 1210
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_RLGYC7  xm7
timestamp 1686918407
transform 1 0 8697 0 1 6561
box -425 -3361 425 3361
use sky130_fd_pr__nfet_01v8_6WGMFU  xm8
timestamp 1686918407
transform 1 0 9655 0 1 3352
box -425 -3352 425 3352
use sky130_fd_pr__res_high_po_0p69_NKSDAM  xR1
timestamp 1686918407
transform 1 0 6235 0 1 4598
box -235 -4598 235 4598
use sky130_fd_pr__res_high_po_0p69_NKSDAM  xR2
timestamp 1686918407
transform 1 0 6599 0 1 4598
box -235 -4598 235 4598
use sky130_fd_pr__res_high_po_0p69_T6SKYN  xR3
timestamp 1686918407
transform 1 0 6963 0 1 4912
box -235 -2598 235 2598
<< labels >>
flabel metal1 6000 -200 6200 0 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 6000 9920 6200 10120 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel via1 9500 10300 9700 10500 0 FreeSans 256 0 0 0 out2
port 4 nsew
flabel via1 7220 -546 7420 -346 0 FreeSans 256 0 0 0 in1
port 2 nsew
flabel via1 8268 -546 8468 -346 0 FreeSans 256 0 0 0 in2
port 3 nsew
<< end >>
