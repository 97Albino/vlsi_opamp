* SPICE3 file created from opamp2.ext - technology: (null)

X0 a_8466_4122# m1_7080_2810.t2 vdd vdd sky130_fd_pr__pfet_01v8
X1 a_8466_4122# in2.t0 m1_7402_2810# gnd sky130_fd_pr__nfet_01v8
X2 vdd m1_7080_2810.t0 m1_7080_2810.t1 vdd sky130_fd_pr__pfet_01v8
R0 in1.n1 in1.t0 30.5835
R1 in1.n1 in1.n0 0.0630003
R2 in1 in1.n1 0.063
R3 m1_7080_2810.n0 m1_7080_2810.t2 257.476
R4 m1_7080_2810.n0 m1_7080_2810.t0 256.43
R5 m1_7080_2810.t1 m1_7080_2810.n0 4.44547
R6 gnd.n24 gnd.n22 1407.97
R7 gnd.n21 gnd.n19 1407.97
R8 gnd.n79 gnd.n71 1054.53
R9 gnd.n98 gnd.n69 1054.53
R10 gnd.n59 gnd.n52 856.876
R11 gnd.n59 gnd.n53 856.876
R12 gnd.n100 gnd.n99 341.692
R13 gnd.n4 gnd.n2 277.202
R14 gnd.n9 gnd.n4 225.369
R15 gnd.n95 gnd.n93 133.363
R16 gnd.n81 gnd.n80 128.221
R17 gnd.n26 gnd.n25 126.942
R18 gnd.n41 gnd.n39 120.094
R19 gnd.n41 gnd.n40 120.094
R20 gnd.n68 gnd.n67 116.6
R21 gnd.n87 gnd.n86 110.629
R22 gnd.n58 gnd.n57 108.808
R23 gnd.n109 gnd.n102 107.203
R24 gnd.n15 gnd.n14 106.564
R25 gnd.n26 gnd.n18 104.99
R26 gnd.n99 gnd.n68 90.673
R27 gnd.n61 gnd.n60 54.8576
R28 gnd.n76 gnd.n75 44.4619
R29 gnd.n6 gnd.n5 39.1337
R30 gnd.n39 gnd.n38 33.8092
R31 gnd.n97 gnd.n96 33.2805
R32 gnd.n96 gnd.n95 33.2805
R33 gnd.n104 gnd.n103 32.1427
R34 gnd.n65 gnd.n64 30.1719
R35 gnd.n80 gnd.n70 27.7338
R36 gnd.n30 gnd.n28 11.9029
R37 gnd.n28 gnd.n15 11.5615
R38 gnd.n11 gnd.n9 9.43605
R39 gnd.n110 gnd.n109 9.3005
R40 gnd.n31 gnd.n30 9.3005
R41 gnd.n63 gnd.n62 9.0005
R42 gnd.n11 gnd.n10 9.0005
R43 gnd.n109 gnd.n108 8.92775
R44 gnd.n49 gnd.n33 8.3605
R45 gnd.n62 gnd.n61 7.8005
R46 gnd.n46 gnd.n43 3.81829
R47 gnd.n49 gnd.n48 3.3605
R48 gnd.n9 gnd.n8 2.8805
R49 gnd.n30 gnd.n29 0.780988
R50 vss gnd.n110 0.492688
R51 gnd.n75 gnd.n72 0.403463
R52 gnd.n110 gnd.n63 0.387219
R53 gnd.n31 gnd.n11 0.284484
R54 gnd.n32 gnd.n31 0.284484
R55 gnd.n93 gnd.n81 0.271878
R56 gnd.n63 gnd.n51 0.114953
R57 gnd.n50 gnd.n32 0.0821406
R58 gnd.n66 gnd.n65 0.079129
R59 gnd.n67 gnd.n66 0.079129
R60 gnd.n75 gnd.n74 0.079129
R61 gnd.n74 gnd.n73 0.079129
R62 gnd.n77 gnd.n76 0.079129
R63 gnd.n78 gnd.n77 0.079129
R64 gnd.n80 gnd.n79 0.079129
R65 gnd.n79 gnd.n78 0.079129
R66 gnd.n98 gnd.n97 0.079129
R67 gnd.n99 gnd.n98 0.079129
R68 gnd.n95 gnd.n94 0.079129
R69 gnd.n81 gnd 0.078625
R70 gnd.n21 gnd.n20 0.0464978
R71 gnd.n25 gnd.n21 0.0464978
R72 gnd.n35 gnd.n34 0.0464978
R73 gnd.n36 gnd.n35 0.0464978
R74 gnd.n24 gnd.n23 0.0464978
R75 gnd.n25 gnd.n24 0.0464978
R76 gnd.n38 gnd.n37 0.0464978
R77 gnd.n37 gnd.n36 0.0464978
R78 gnd.n108 gnd.n107 0.0464978
R79 gnd.n107 gnd.n106 0.0464978
R80 gnd.n105 gnd.n104 0.0464978
R81 gnd.n106 gnd.n105 0.0464978
R82 gnd.n51 gnd.n50 0.0333125
R83 gnd.n42 gnd.n41 0.0286765
R84 gnd.n43 gnd.n42 0.0286765
R85 gnd.n56 gnd.n55 0.0286765
R86 gnd.n57 gnd.n56 0.0286765
R87 gnd.n17 gnd.n16 0.0286765
R88 gnd.n18 gnd.n17 0.0286765
R89 gnd.n7 gnd.n6 0.0250974
R90 gnd.n2 gnd.n1 0.0250016
R91 gnd.n1 gnd.n0 0.0250016
R92 gnd.n48 gnd.n47 0.0250016
R93 gnd.n47 gnd.n46 0.0250016
R94 gnd.n8 gnd.n7 0.0250016
R95 gnd.n45 gnd.n44 0.0250016
R96 gnd.n46 gnd.n45 0.0250016
R97 gnd.n59 gnd.n54 0.00687366
R98 gnd.n59 gnd.n58 0.00687366
R99 gnd.n102 gnd.n101 0.00687366
R100 gnd.n101 gnd.n100 0.00687366
R101 gnd.n28 gnd.n27 0.00687366
R102 gnd.n27 gnd.n26 0.00687366
R103 gnd.n60 gnd.n59 0.00368683
R104 gnd.n86 gnd.n85 0.00326136
R105 gnd.n85 gnd.n84 0.00326136
R106 gnd.n83 gnd.n82 0.00326136
R107 gnd.n84 gnd.n83 0.00326136
R108 gnd.n4 gnd.n3 0.00261132
R109 gnd.n14 gnd.n13 0.00261132
R110 gnd.n13 gnd.n12 0.00261132
R111 gnd.n88 gnd.n87 0.00202003
R112 gnd.n91 gnd.n88 0.00202003
R113 gnd.n90 gnd.n89 0.00202003
R114 gnd.n91 gnd.n90 0.00202003
R115 gnd.n93 gnd.n92 0.00202003
R116 gnd.n92 gnd.n91 0.00202003
R117 gnd.n50 gnd.n49 0.000500017
R118 in2.n1 in2.t0 30.5858
R119 in2.n1 in2.n0 0.0630003
R120 in2 in2.n1 0.063
R121 vdd.n22 vdd.n20 857.648
R122 vdd.n8 vdd.n2 857.648
R123 vdd.n18 vdd.n11 108.251
R124 vdd.n19 vdd.n18 105.052
R125 vdd.n10 vdd.n9 44.4348
R126 vdd.n11 vdd.n10 41.3262
R127 vdd.n31 vdd.n30 38.4785
R128 vdd.n31 vdd.n1 14.2005
R129 vdd.n30 vdd.n24 10.8827
R130 vdd vdd.n31 1.02667
R131 vdd.n24 vdd.n19 0.190047
R132 vdd.n10 vdd.n8 0.0150463
R133 vdd.n8 vdd.n7 0.0150463
R134 vdd.n7 vdd.n4 0.0150463
R135 vdd.n4 vdd.n3 0.0150463
R136 vdd.n24 vdd.n22 0.0150463
R137 vdd.n22 vdd.n21 0.0150463
R138 vdd.n24 vdd.n23 0.0150463
R139 vdd.n6 vdd.n5 0.00824837
R140 vdd.n7 vdd.n6 0.00824837
R141 vdd.n1 vdd.n0 0.00824837
R142 vdd.n13 vdd.n12 0.00249866
R143 vdd.n16 vdd.n13 0.00249866
R144 vdd.n18 vdd.n17 0.00249866
R145 vdd.n17 vdd.n16 0.00249866
R146 vdd.n15 vdd.n14 0.00249866
R147 vdd.n16 vdd.n15 0.00249866
R148 vdd.n29 vdd.n28 0.00159127
R149 vdd.n26 vdd.n25 0.00116581
R150 vdd.n27 vdd.n26 0.00116581
R151 vdd.n30 vdd.n29 0.00116581
R152 vdd.n28 vdd.n27 0.00107455
R153 out2 out2.n0 0.1255
C0 out2.n0 0 0.115f **FLOATING
C1 out2 0 16.1f **FLOATING
C2 vdd.n0 0 1.62f **FLOATING
C3 vdd.n1 0 0.874f **FLOATING
C4 vdd.n2 0 0.0132f **FLOATING
C5 vdd.n3 0 0.0283f **FLOATING
C6 vdd.n4 0 0.0134f **FLOATING
C7 vdd.n5 0 0.0698f **FLOATING
C8 vdd.n6 0 0.0595f **FLOATING
C9 vdd.n7 0 0.581f **FLOATING
C10 vdd.n8 0 0.0134f **FLOATING
C11 vdd.n9 0 0.0173f **FLOATING
C12 vdd.n10 0 0.00777f **FLOATING
C13 vdd.n11 0 0.0512f **FLOATING
C14 vdd.n12 0 0.0426f **FLOATING
C15 vdd.n13 0 0.0225f **FLOATING
C16 vdd.n14 0 0.0185f **FLOATING
C17 vdd.n15 0 0.0185f **FLOATING
C18 vdd.n16 0 1.06f **FLOATING
C19 vdd.n17 0 0.0225f **FLOATING
C20 vdd.n18 0 0.0773f **FLOATING
C21 vdd.n19 0 0.071f **FLOATING
C22 vdd.n20 0 0.0132f **FLOATING
C23 vdd.n21 0 0.978f **FLOATING
C24 vdd.n22 0 0.0134f **FLOATING
C25 vdd.n23 0 0.0134f **FLOATING
C26 vdd.n24 0 0.27f **FLOATING
C27 vdd.n25 0 1.64f **FLOATING
C28 vdd.n26 0 0.059f **FLOATING
C29 vdd.n27 0 1.96f **FLOATING
C30 vdd.n29 0 0.059f **FLOATING
C31 vdd.n30 0 1.16f **FLOATING
C32 vdd.n31 0 2.9f **FLOATING
C33 vdd 0 0.354f **FLOATING
C34 m1_7080_2810.t2 0 0.589f **FLOATING
C35 m1_7080_2810.t0 0 0.588f **FLOATING
C36 m1_7080_2810.n0 0 1.15f **FLOATING
C37 m1_7080_2810.t1 0 0.275f **FLOATING
