magic
tech sky130B
magscale 1 2
timestamp 1685704482
<< checkpaint >>
rect 8204 7203 11194 11256
rect 7887 3540 11194 7203
rect -1260 -3260 1460 1460
rect 7887 -513 10877 3540
<< nwell >>
rect 10200 7038 12050 11322
rect 11200 4840 12050 7038
rect 10802 4794 12050 4840
rect 11200 4600 12050 4794
<< pwell >>
rect 11134 3200 11194 3632
rect 11060 3140 11194 3200
<< locali >>
rect 8160 11480 13660 11520
rect 8160 11280 8500 11480
rect 13560 11280 13660 11480
rect 8160 11240 13660 11280
rect 8160 10400 11480 11240
rect 8160 9920 9934 10034
rect 8160 900 8446 9920
rect 8760 900 8820 9920
rect 9120 4880 9540 9920
rect 9860 4880 9934 9920
rect 9120 4600 9934 4880
rect 10200 6960 11480 10400
rect 10200 4680 10280 6960
rect 11208 4680 11480 6960
rect 12180 7600 13660 11240
rect 12180 4680 12320 7600
rect 10200 4600 12320 4680
rect 12560 7260 13660 7304
rect 9120 900 9200 4600
rect 12560 4300 12680 7260
rect 8160 800 9200 900
rect 9420 4120 12680 4300
rect 9420 3500 10280 4120
rect 10700 3500 10780 4120
rect 11200 3500 12680 4120
rect 9420 2950 12680 3500
rect 9420 680 9500 2950
rect 9920 680 10400 2950
rect 11080 680 12680 2950
rect 13360 680 13660 7260
rect 8160 640 13660 680
rect 8160 440 8500 640
rect 13540 440 13660 640
rect 8160 400 13660 440
<< viali >>
rect 8500 11280 13560 11480
rect 8500 440 13540 640
<< metal1 >>
rect 8160 11480 13660 11520
rect 8160 11280 8500 11480
rect 13560 11280 13660 11480
rect 8160 11252 11780 11280
rect 11860 11252 13660 11280
rect 8160 11240 13660 11252
rect 8532 9398 8670 11240
rect 8896 9398 9768 9830
rect 10280 6820 10338 11240
rect 8160 5530 8400 5890
rect 9620 4966 9630 5398
rect 9768 4966 9778 5398
rect 10280 4818 10390 6820
rect 10456 4778 10536 6860
rect 10602 6818 10720 6820
rect 10648 4822 10720 6818
rect 10602 4800 10720 4822
rect 10790 4940 10876 6820
rect 10790 4880 10800 4940
rect 10860 4880 10876 4940
rect 10790 4818 10876 4880
rect 10602 4778 10620 4800
rect 10400 4740 10620 4778
rect 10680 4778 10720 4800
rect 10940 4778 11020 6860
rect 11140 6820 11206 11240
rect 11520 11042 11530 11102
rect 11590 11042 11600 11102
rect 11086 4818 11206 6820
rect 11630 4778 11728 11144
rect 11774 5820 11784 6140
rect 11864 5820 11874 6140
rect 11920 4778 12018 11144
rect 12050 11042 12060 11102
rect 12120 11042 12130 11102
rect 10680 4740 11078 4778
rect 10400 4732 11078 4740
rect 11600 4732 12050 4778
rect 10284 3200 10344 3692
rect 10454 3600 10534 4060
rect 10602 3880 10690 3990
rect 10648 3840 10690 3880
rect 10610 3780 10620 3840
rect 10680 3780 10690 3840
rect 10648 3740 10690 3780
rect 10602 3632 10690 3740
rect 10790 3840 10830 3990
rect 10790 3780 10800 3840
rect 10860 3780 10870 3840
rect 10790 3632 10830 3780
rect 10942 3600 11022 4062
rect 10398 3536 10408 3600
rect 10584 3536 10594 3600
rect 10884 3536 10894 3600
rect 11070 3536 11080 3600
rect 11134 3200 11194 3692
rect 10284 3140 11194 3200
rect 9656 2842 9666 2922
rect 9746 2842 9756 2922
rect 9508 2730 9518 2810
rect 9598 2730 9608 2810
rect 8532 966 9034 1398
rect 9656 778 9754 2842
rect 10284 2810 10344 3140
rect 10520 2922 10970 2940
rect 10520 2908 10706 2922
rect 10520 2842 10574 2908
rect 10564 2828 10574 2842
rect 10654 2842 10706 2908
rect 10786 2908 10970 2922
rect 10786 2844 10854 2908
rect 10786 2842 10830 2844
rect 10844 2842 10854 2844
rect 10654 2828 10664 2842
rect 9852 860 9914 2810
rect 10284 2750 10466 2810
rect 9810 810 9914 860
rect 9862 680 9914 810
rect 10564 778 10664 2828
rect 10840 2828 10854 2842
rect 10934 2842 10970 2908
rect 10934 2828 10946 2842
rect 10696 840 10706 916
rect 10786 840 10796 916
rect 10840 778 10946 2828
rect 11134 2810 11194 3140
rect 11026 2750 11194 2810
rect 12720 810 12730 870
rect 12790 810 12800 870
rect 12840 780 12940 7126
rect 12974 5820 12984 6140
rect 13064 5820 13074 6140
rect 13120 780 13220 7126
rect 13430 5880 13440 6080
rect 13640 5880 13650 6080
rect 13250 810 13260 870
rect 13320 810 13330 870
rect 10564 772 10598 778
rect 10820 776 10830 778
rect 12796 722 12994 780
rect 12984 720 12994 722
rect 13054 722 13254 780
rect 13054 720 13064 722
rect 8160 670 13660 680
rect 8160 640 10706 670
rect 10786 660 13660 670
rect 10786 640 12980 660
rect 13060 640 13660 660
rect 8160 440 8500 640
rect 13540 440 13660 640
rect 8160 400 13660 440
rect 0 0 200 200
rect 10386 100 10396 300
rect 10596 100 10606 300
rect 10874 90 10884 290
rect 11084 90 11094 290
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
<< via1 >>
rect 11780 11280 11860 11332
rect 11780 11252 11860 11280
rect 9630 4966 9768 5398
rect 10800 4880 10860 4940
rect 10620 4740 10680 4800
rect 11530 11042 11590 11102
rect 11784 5820 11864 6140
rect 12060 11042 12120 11102
rect 10620 3780 10680 3840
rect 10800 3780 10860 3840
rect 10408 3536 10584 3600
rect 10894 3536 11070 3600
rect 9666 2842 9746 2922
rect 9518 2730 9598 2810
rect 10574 2828 10654 2908
rect 10706 2842 10786 2922
rect 10854 2828 10934 2908
rect 10706 840 10786 916
rect 12730 810 12790 870
rect 12984 5820 13064 6140
rect 13440 5880 13640 6080
rect 13260 810 13320 870
rect 12994 720 13054 780
rect 10706 640 10786 670
rect 12980 640 13060 660
rect 10706 594 10786 640
rect 12980 580 13060 640
rect 10396 100 10596 300
rect 10884 90 11084 290
<< metal2 >>
rect 11780 11332 11860 11342
rect 11780 11242 11860 11252
rect 11530 11102 11590 11112
rect 11530 11032 11590 11042
rect 12060 11102 12120 11112
rect 12060 11032 12120 11042
rect 11784 6140 13660 6150
rect 11864 5820 12984 6140
rect 13064 6080 13660 6140
rect 13064 5880 13440 6080
rect 13640 5880 13660 6080
rect 13064 5820 13660 5880
rect 11784 5810 13660 5820
rect 9630 5398 9768 5408
rect 9518 4966 9630 5398
rect 9768 4966 9840 5398
rect 9518 2932 9840 4966
rect 10800 4940 10860 4950
rect 10620 4800 10680 4810
rect 10620 3840 10680 4740
rect 10620 3770 10680 3780
rect 10800 4784 10860 4880
rect 10800 3840 10860 4724
rect 11794 4786 11854 4796
rect 11794 4716 11854 4726
rect 10800 3770 10860 3780
rect 10408 3600 10584 3610
rect 10408 3526 10584 3536
rect 10894 3600 11070 3610
rect 10894 3526 11070 3536
rect 9518 2922 13120 2932
rect 9518 2842 9666 2922
rect 9746 2908 10706 2922
rect 9746 2842 10574 2908
rect 9518 2828 10574 2842
rect 10654 2842 10706 2908
rect 10786 2908 13120 2922
rect 10786 2842 10854 2908
rect 10654 2828 10854 2842
rect 10934 2828 13120 2908
rect 9518 2810 13120 2828
rect 9598 2730 13120 2810
rect 9518 2720 13120 2730
rect 10706 916 10786 926
rect 10706 670 10786 840
rect 12730 870 12790 880
rect 12730 800 12790 810
rect 12940 780 13120 2720
rect 13260 870 13320 880
rect 13260 800 13320 810
rect 12940 720 12994 780
rect 13054 720 13120 780
rect 12940 710 13120 720
rect 10706 584 10786 594
rect 12980 660 13060 670
rect 12980 570 13060 580
rect 10396 300 10596 310
rect 10396 90 10596 100
rect 10884 290 11084 300
rect 10884 80 11084 90
<< via2 >>
rect 11780 11252 11860 11332
rect 11530 11042 11590 11102
rect 12060 11042 12120 11102
rect 10800 4724 10860 4784
rect 11794 4726 11854 4786
rect 10408 3536 10582 3600
rect 10894 3536 11070 3600
rect 12730 810 12790 870
rect 13260 810 13320 870
rect 12980 580 13060 660
rect 10396 100 10594 300
rect 10884 90 11084 290
<< metal3 >>
rect 11770 11332 11870 11337
rect 11770 11252 11780 11332
rect 11860 11252 11870 11332
rect 11770 11247 11870 11252
rect 11780 11108 11860 11247
rect 11520 11102 12130 11108
rect 11520 11042 11530 11102
rect 11590 11042 12060 11102
rect 12120 11042 12130 11102
rect 11520 11036 12130 11042
rect 10780 4786 11880 4800
rect 10780 4784 11794 4786
rect 10780 4724 10800 4784
rect 10860 4726 11794 4784
rect 11854 4726 11880 4786
rect 10860 4724 11880 4726
rect 10780 4700 11880 4724
rect 10384 3600 10604 3606
rect 10384 3536 10408 3600
rect 10582 3536 10604 3600
rect 10884 3600 11080 3605
rect 10884 3596 10894 3600
rect 10384 300 10604 3536
rect 10384 100 10396 300
rect 10594 100 10604 300
rect 10384 95 10604 100
rect 10874 3536 10894 3596
rect 11070 3596 11080 3600
rect 11070 3536 11094 3596
rect 10874 290 11094 3536
rect 12720 870 13330 880
rect 12720 810 12730 870
rect 12790 810 13260 870
rect 13320 810 13330 870
rect 12720 800 13330 810
rect 12980 665 13060 800
rect 12970 660 13070 665
rect 12970 580 12980 660
rect 13060 580 13070 660
rect 12970 575 13070 580
rect 10874 90 10884 290
rect 11084 90 11094 290
rect 10874 85 11094 90
use sky130_fd_pr__res_high_po_0p69_YVB7ZU  sky130_fd_pr__res_high_po_0p69_YVB7ZU_0
timestamp 1683799460
transform 1 0 9699 0 1 7398
box -235 -2598 235 2598
use sky130_fd_pr__nfet_01v8_34YWRA  xm1
timestamp 1683799460
transform 1 0 10496 0 1 3811
box -296 -389 296 389
use sky130_fd_pr__nfet_01v8_34YWRA  xm2
timestamp 1683799460
transform 1 0 10982 0 1 3811
box -296 -389 296 389
use sky130_fd_pr__pfet_01v8_GGAEPD  xm3
timestamp 1683799460
transform 1 0 10496 0 1 5819
box -296 -1219 296 1219
use sky130_fd_pr__pfet_01v8_GGAEPD  xm4
timestamp 1683799460
transform 1 0 10982 0 1 5819
box -296 -1219 296 1219
use sky130_fd_pr__nfet_01v8_EF4BLE  xm5
timestamp 1683799460
transform -1 0 10745 0 -1 1810
box -425 -1210 425 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  xm6
timestamp 1683799460
transform -1 0 9704 0 -1 1810
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_RLGYC7  xm7
timestamp 1683799460
transform -1 0 11825 0 -1 7961
box -425 -3361 425 3361
use sky130_fd_pr__nfet_01v8_6WGMFU  xm8
timestamp 1683799460
transform -1 0 13025 0 -1 3952
box -425 -3352 425 3352
use sky130_fd_pr__res_high_po_0p69_NKSDAM  xR1
timestamp 1683799460
transform 1 0 8601 0 1 5398
box -235 -4598 235 4598
use sky130_fd_pr__res_high_po_0p69_NKSDAM  xR2
timestamp 1683799460
transform 1 0 8965 0 1 5398
box -235 -4598 235 4598
use sky130_fd_pr__res_high_po_0p69_YVB7ZU  xR3
timestamp 1683799460
transform 1 0 9382 0 1 3345
box -235 -2598 235 2598
<< labels >>
flabel metal1 8240 11280 8440 11480 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel via1 10884 90 11084 290 0 FreeSans 256 0 0 0 in2
port 3 nsew
flabel via1 10396 100 10596 300 0 FreeSans 256 0 0 0 in1
port 2 nsew
flabel via1 13440 5880 13640 6080 0 FreeSans 256 0 0 0 out2
port 4 nsew
flabel metal1 8180 5610 8380 5810 0 FreeSans 256 0 0 0 gnd
flabel metal1 8240 440 8440 640 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 vdd
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 vss
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 gnd
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 in1
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 in2
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 out2
port 5 nsew
<< end >>
