magic
tech sky130B
magscale 1 2
timestamp 1683799460
<< pwell >>
rect -296 -389 296 389
<< nmos >>
rect -100 -179 100 179
<< ndiff >>
rect -158 167 -100 179
rect -158 -167 -146 167
rect -112 -167 -100 167
rect -158 -179 -100 -167
rect 100 167 158 179
rect 100 -167 112 167
rect 146 -167 158 167
rect 100 -179 158 -167
<< ndiffc >>
rect -146 -167 -112 167
rect 112 -167 146 167
<< psubdiff >>
rect -260 319 -164 353
rect 164 319 260 353
rect -260 257 -226 319
rect 226 257 260 319
rect -260 -319 -226 -257
rect 226 -319 260 -257
rect -260 -353 -164 -319
rect 164 -353 260 -319
<< psubdiffcont >>
rect -164 319 164 353
rect -260 -257 -226 257
rect 226 -257 260 257
rect -164 -353 164 -319
<< poly >>
rect -100 251 100 267
rect -100 217 -84 251
rect 84 217 100 251
rect -100 179 100 217
rect -100 -217 100 -179
rect -100 -251 -84 -217
rect 84 -251 100 -217
rect -100 -267 100 -251
<< polycont >>
rect -84 217 84 251
rect -84 -251 84 -217
<< locali >>
rect -260 319 -164 353
rect 164 319 260 353
rect -260 257 -226 319
rect 226 257 260 319
rect -100 217 -84 251
rect 84 217 100 251
rect -146 167 -112 183
rect -146 -183 -112 -167
rect 112 167 146 183
rect 112 -183 146 -167
rect -100 -251 -84 -217
rect 84 -251 100 -217
rect -260 -319 -226 -257
rect 226 -319 260 -257
rect -260 -353 -164 -319
rect 164 -353 260 -319
<< viali >>
rect -84 217 84 251
rect -146 -167 -112 167
rect 112 -167 146 167
rect -84 -251 84 -217
<< metal1 >>
rect -96 251 96 257
rect -96 217 -84 251
rect 84 217 96 251
rect -96 211 96 217
rect -152 167 -106 179
rect -152 -167 -146 167
rect -112 -167 -106 167
rect -152 -179 -106 -167
rect 106 167 152 179
rect 106 -167 112 167
rect 146 -167 152 167
rect 106 -179 152 -167
rect -96 -217 96 -211
rect -96 -251 -84 -217
rect 84 -251 96 -217
rect -96 -257 96 -251
<< properties >>
string FIXED_BBOX -243 -336 243 336
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.79 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
