* SPICE3 file created from opamp.ext - technology: sky130B

.subckt opamp vdd vss in1 in2 out2
X0 a_8668_3322# in2 m1_7702_2524# vss sky130_fd_pr__nfet_01v8 ad=0.519 pd=4.16 as=0.519 ps=4.16 w=1.79 l=1
X1 vdd m1_8030_3374# m1_8030_3374# vdd sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.6 as=2.9 ps=20.6 w=10 l=1
X2 a_8668_3322# m1_8030_3374# vdd vdd sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.6 as=2.9 ps=20.6 w=10 l=1
X3 m1_7702_2524# m1_6894_2242# vss vss sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.3 as=2.9 ps=20.6 w=10 l=1
X4 vss m1_6894_2242# m1_7702_2524# vss sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.6 as=1.45 ps=10.3 w=10 l=1
X5 m1_6894_2242# m1_6894_2242# vss vss sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.6 as=2.9 ps=20.6 w=10 l=1
X6 vdd a_8668_3322# out2 vdd sky130_fd_pr__pfet_01v8 ad=9.11 pd=63.4 as=4.56 ps=31.7 w=31.4 l=1
X7 out2 a_8668_3322# vdd vdd sky130_fd_pr__pfet_01v8 ad=4.56 pd=31.7 as=9.11 ps=63.4 w=31.4 l=1
X8 out2 m1_6894_2242# vss vss sky130_fd_pr__nfet_01v8 ad=4.56 pd=31.7 as=9.11 ps=63.4 w=31.4 l=1
X9 vss m1_6894_2242# out2 vss sky130_fd_pr__nfet_01v8 ad=9.11 pd=63.4 as=4.56 ps=31.7 w=31.4 l=1
X10 m1_7702_2524# in1 m1_8030_3374# vss sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.79 l=1
X11 m1_6166_166# m1_6530_8598# vss sky130_fd_pr__res_high_po_0p69 l=40
X12 m1_6166_166# vdd vss sky130_fd_pr__res_high_po_0p69 l=40
X13 m1_6894_2242# m1_6530_8598# vss sky130_fd_pr__res_high_po_0p69 l=20
.ends
